module DSP(A,B,D,C,CLK,CARRYIN,OPMODE,BCIN,RSTA,RSTB,RSTM,RSTP,RSTC,RSTD,RSTCARRYIN,RSTOPMODE,CEA,CEB,CEM,CEP,CEC,CED,CECARRYIN,CEOPMODE,PCIN,
                BCOUT,PCOUT,P,M,CARRYOUT,CARRYOUTF);

input [17:0] A,B,D,BCIN;
input [47:0] C , PCIN;
input [7:0]  OPMODE;
input CARRYIN,CLK,RSTA,RSTB,RSTM,RSTP,RSTC,RSTD,RSTCARRYIN,RSTOPMODE,CEA,CEB,CEM,CEP,CEC,CED,CECARRYIN,CEOPMODE ;
output [17:0] BCOUT;
output  [35:0] M;
output  [47:0] P ,PCOUT;
output  CARRYOUT,CARRYOUTF;

parameter RSTTYPE = "SYNC";

generate 
    if( RSTTYPE == "SYNC")
      DSP_sync DSPS(A,B,D,C,CLK,CARRYIN,OPMODE,BCIN,RSTA,RSTB,RSTM,RSTP,RSTC,RSTD,RSTCARRYIN,RSTOPMODE,CEA,CEB,CEM,CEP,CEC,CED,CECARRYIN,CEOPMODE,PCIN,
                BCOUT,PCOUT,P,M,CARRYOUT,CARRYOUTF);
   else 
      DSP_async DSPA(A,B,D,C,CLK,CARRYIN,OPMODE,BCIN,RSTA,RSTB,RSTM,RSTP,RSTC,RSTD,RSTCARRYIN,RSTOPMODE,CEA,CEB,CEM,CEP,CEC,CED,CECARRYIN,CEOPMODE,PCIN,
                BCOUT,PCOUT,P,M,CARRYOUT,CARRYOUTF);
endgenerate

endmodule



